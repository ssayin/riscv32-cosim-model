module riscv_core_wrapper ();

  // riscv_core riscv_core_0 (
  // .clk          (clk_100MHz),
  // .rst_n        (reset_rtl_0),
  // .axi_arddr_f  (S_AXI_araddr),
  // .axi_arburst_f(S_AXI_arburst),
  // .axi_arcache_f(S_AXI_arcache),
  // .axi_arlen_f  (S_AXI_arlen),
  // .axi_arlock_f (S_AXI_arlock),
  // .axi_arprot_f (S_AXI_arprot),
  // .axi_arready_f(S_AXI_arready),
  // .axi_arsize_f (S_AXI_arsize),
  // .axi_arvalid_f(S_AXI_arvalid),
  // .axi_awaddr_f (S_AXI_awaddr),
  // .axi_awburst_f(S_AXI_awburst),
  // .axi_awcache_f(S_AXI_awcache),
  // .axi_awlen_f  (S_AXI_awlen),
  // .axi_awlock_f (S_AXI_awlock),
  // .axi_awprot_f (S_AXI_awprot),
  // .axi_awready_f(S_AXI_awready),
  // .axi_awsize_f (S_AXI_awsize),
  // .axi_awvalid_f(S_AXI_awvalid),
  // .axi_bready_f (S_AXI_bready),
  // .axi_bresp_f  (S_AXI_bresp),
  // .axi_bvalid_f (S_AXI_bvalid),
  // .axi_rdata_f  (S_AXI_rdata),
  // .axi_rlast_f  (S_AXI_rlast),
  // .axi_rready_f (S_AXI_rready),
  // .axi_rresp_f  (S_AXI_rresp),
  // .axi_rvalid_f (S_AXI_rvalid),
  // .axi_wdata_f  (S_AXI_wdata),
  // .axi_wlast_f  (S_AXI_wlast),
  // .axi_wready_f (S_AXI_wready),
  // .axi_wstrb_f  (S_AXI_wstrb),
  // .axi_wvalid_f (S_AXI_wvalid)
  // );

endmodule

