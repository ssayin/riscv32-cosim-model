// SPDX-FileCopyrightText: 2023 Serdar Sayın <https://serdarsayin.com>
//
// SPDX-License-Identifier: Apache-2.0

//=============================================================================
// Project  : src/tb/uvm_bfm
//
// File Name: axi4ar_sequencer.sv
//
// Author   : Name   : Serdar Sayın
//            Email  : serdarsayin@pm.me
//            Year   : 2023
//
// Version:   0.1
//
// Code created by Easier UVM Code Generator version 2017-01-19 on Mon Aug 14 04:22:47 2023
//=============================================================================
// Description: Sequencer for axi4ar
//=============================================================================

`ifndef AXI4AR_SEQUENCER_SV
`define AXI4AR_SEQUENCER_SV

// Sequencer class is specialization of uvm_sequencer
typedef uvm_sequencer #(axi4ar_tx) axi4ar_sequencer_t;


`endif // AXI4AR_SEQUENCER_SV

