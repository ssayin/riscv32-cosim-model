// SPDX-FileCopyrightText: 2023 Serdar Sayın <https://serdarsayin.com>
//
// SPDX-License-Identifier: Apache-2.0

//=============================================================================
// Project  : src/tb/uvm_top
//
// File Name: _if.sv
//
// Author   : Name   : Serdar Sayın
//            Email  : serdarsayin@pm.me
//            Year   : 2023
//
// Version:   0.1
//
// Code created by Easier UVM Code Generator version 2017-01-19 on Sat Aug 12 02:59:40 2023
//=============================================================================
// Description: Signal interface for agent 
//=============================================================================

`ifndef _IF_SV
`define _IF_SV

interface (); 

  timeunit      1ns;
  timeprecision 1ps;

  import _pkg::*;


  // You can insert properties and assertions here

endinterface : 

`endif // _IF_SV

