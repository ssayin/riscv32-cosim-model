// SPDX-FileCopyrightText: 2023 Serdar Sayın <https://serdarsayin.com>
//
// SPDX-License-Identifier: Apache-2.0

//=============================================================================
// Project  : src/tb/uvm_top
//
// File Name: riscv_core_sequencer.sv
//
// Author   : Name   : Serdar Sayın
//            Email  : serdarsayin@pm.me
//            Year   : 2023
//
// Version:   0.1
//
// Code created by Easier UVM Code Generator version 2017-01-19 on Sat Aug 12 03:33:22 2023
//=============================================================================
// Description: Sequencer for riscv_core
//=============================================================================

`ifndef RISCV_CORE_SEQUENCER_SV
`define RISCV_CORE_SEQUENCER_SV

// Sequencer class is specialization of uvm_sequencer
typedef uvm_sequencer #(riscv_core_tx) riscv_core_sequencer_t;


`endif // RISCV_CORE_SEQUENCER_SV

