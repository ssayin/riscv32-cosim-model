// SPDX-FileCopyrightText: 2023 Serdar Sayın <https://serdarsayin.com>
//
// SPDX-License-Identifier: Apache-2.0

// TODO: what are trade-off btw. decompress expansion
// VS decode right justified w/ comp switch?
module ifu_aln ();
endmodule
