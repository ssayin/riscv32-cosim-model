module top_level ();

endmodule
