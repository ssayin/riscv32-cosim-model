// SPDX-FileCopyrightText: 2023 Serdar Sayın <https://serdarsayin.com>
//
// SPDX-License-Identifier: Apache-2.0

//=============================================================================
// Project  : ../tb/uvm_top
//
// File Name: top_config.sv
//
// Author   : Name   : Serdar Sayın
//            Email  : serdarsayin@pm.me
//            Year   : 2023
//
// Version:   0.1
//
// Code created by Easier UVM Code Generator version 2017-01-19 on Wed Aug  2 13:55:59 2023
//=============================================================================
// Description: Configuration for top
//=============================================================================

`ifndef TOP_CONFIG_SV
`define TOP_CONFIG_SV

// You can insert code here by setting top_env_config_inc_before_class in file common.tpl

class top_config extends uvm_object;

  // Do not register config class with the factory

  rand axi4master_config  m_axi4master_0_config;
  rand axi4master_config  m_axi4master_1_config;

  // You can insert variables here by setting config_var in file common.tpl

  // You can remove new by setting top_env_config_generate_methods_inside_class = no in file common.tpl

  extern function new(string name = "");

  // You can insert code here by setting top_env_config_inc_inside_class in file common.tpl

endclass : top_config 


// You can remove new by setting top_env_config_generate_methods_after_class = no in file common.tpl

function top_config::new(string name = "");
  super.new(name);

  m_axi4master_0_config                 = new("m_axi4master_0_config");
  m_axi4master_0_config.is_active       = UVM_ACTIVE;                  
  m_axi4master_0_config.checks_enable   = 1;                           
  m_axi4master_0_config.coverage_enable = 1;                           

  m_axi4master_1_config                 = new("m_axi4master_1_config");
  m_axi4master_1_config.is_active       = UVM_ACTIVE;                  
  m_axi4master_1_config.checks_enable   = 1;                           
  m_axi4master_1_config.coverage_enable = 1;                           

  // You can insert code here by setting top_env_config_append_to_new in file common.tpl

endfunction : new


// You can insert code here by setting top_env_config_inc_after_class in file common.tpl

`endif // TOP_CONFIG_SV

