module fpga_top (
  input logic clk,
  input logic rst_n
);

endmodule
