`ifndef DEC_DECODE_TEST_LIST
`define DEC_DECODE_TEST_LIST

package dec_decode_test_list;

  import uvm_pkg::*;
  `include "uvm_macros.svh"

  import dec_decode_env_pkg::*;
  import dec_decode_seq_list::*;

  `include "dec_decode_basic_test.sv"
  `include "dec_decode_from_file_test.sv"

endpackage : dec_decode_test_list

`endif



