../../../../src/rtl/include/riscv_opcodes.svh