  riscv_core_ref_model  m_ref_model;
  riscv_core_scoreboard m_scoreboard;

  // riscv_core_coverage #(riscv_core_transaction) coverage;
