module tb_top_level;

  logic clk;
  logic rst_n;

  top_level top_level_0 (.*);

endmodule
