// SPDX-FileCopyrightText: 2023 Serdar Sayın <https://serdarsayin.com>
//
// SPDX-License-Identifier: Apache-2.0

module axi2apb #(
    parameter int ID       = 1,
    parameter int AXI_ADDR = 32,
    parameter int AXI_DATA = 32,
    parameter int APB_ADDR = 32,
    parameter int APB_DATA = 32
) (
  input  logic       clk,
  input  logic       rst_n,
  output logic       awready,
  output logic       bvalid,
  output logic       bid,
  output logic [1:0] bresp,
  output logic       arready,
  output logic       rvalid,
  output logic       rid,
  output logic       rdata,
  output logic [1:0] rresp,
  output logic       rlast,
  output logic       paddr,
  output logic [2:0] prot,
  output logic       penable,
  output logic       pwrite,
  output logic       pwdata,
  output logic [1:0] pstrb,
  output logic       psel,
  input  logic       awvalid,
  input  logic       awid,
  input  logic       awaddr,
  input  logic [7:0] awlen,
  input  logic [2:0] awsize,
  input  logic [1:0] awburst,
  input  logic       awlock,
  input  logic [3:0] awcache,
  input  logic [2:0] awprot,
  input  logic [3:0] awqos,
  input  logic [3:0] awregion,
  input  logic       wvalid,
  input  logic       wdata,
  input  logic [3:0] wstrb,
  input  logic       wlast,
  input  logic       bready,
  input  logic       arvalid,
  input  logic       arid,
  input  logic       araddr,
  input  logic [7:0] arlen,
  input  logic [2:0] arsize,
  input  logic [1:0] arburst,
  input  logic       arlock,
  input  logic [3:0] arcache,
  input  logic [2:0] arprot,
  input  logic [3:0] arqos,
  input  logic [3:0] arregion,
  input  logic       rready,
  input  logic       pready,
  input  logic       prdata,
  input  logic       pslverr
);

endmodule
