// SPDX-FileCopyrightText: 2023 Serdar Sayın <https://serdarsayin.com>
//
// SPDX-License-Identifier: Apache-2.0

package wb_stage_pkg;

  import uvm_pkg::*;

  `include "uvm_macros.svh"

  `include "wb_stage_agent.sv"
  `include "wb_stage_monitor.sv"
  `include "wb_stage_driver.sv"
  `include "wb_stage_sequencer.sv"
  `include "wb_stage_sequence.sv"

endpackage : wb_stage_pkg
