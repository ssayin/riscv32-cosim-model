tb_dec_decode.sv