// SPDX-FileCopyrightText: 2023 Serdar Sayın <https://serdarsayin.com>
//
// SPDX-License-Identifier: Apache-2.0

//=============================================================================
// Project  : src/tb/uvm_top
//
// File Name: _sequencer.sv
//
// Author   : Name   : Serdar Sayın
//            Email  : serdarsayin@pm.me
//            Year   : 2023
//
// Version:   0.1
//
// Code created by Easier UVM Code Generator version 2017-01-19 on Sat Aug 12 02:59:40 2023
//=============================================================================
// Description: Sequencer for 
//=============================================================================

`ifndef _SEQUENCER_SV
`define _SEQUENCER_SV

// Sequencer class is specialization of uvm_sequencer
typedef uvm_sequencer #() _sequencer_t;


`endif // _SEQUENCER_SV

