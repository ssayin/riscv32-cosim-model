// SPDX-FileCopyrightText: 2023 Serdar Sayın <https://serdarsayin.com>
//
// SPDX-License-Identifier: Apache-2.0

package defs_pkg;

  // verilog_format: off
  parameter logic [31:0] ADD        = 32'b0000000??????????000?????0110011;
  parameter logic [31:0] ADDI       = 32'b?????????????????000?????0010011;
  parameter logic [31:0] AND        = 32'b0000000??????????111?????0110011;
  parameter logic [31:0] ANDI       = 32'b?????????????????111?????0010011;
  parameter logic [31:0] AUIPC      = 32'b?????????????????????????0010111;
  parameter logic [31:0] BEQ        = 32'b?????????????????000?????1100011;
  parameter logic [31:0] BGE        = 32'b?????????????????101?????1100011;
  parameter logic [31:0] BGEU       = 32'b?????????????????111?????1100011;
  parameter logic [31:0] BLT        = 32'b?????????????????100?????1100011;
  parameter logic [31:0] BLTU       = 32'b?????????????????110?????1100011;
  parameter logic [31:0] BNE        = 32'b?????????????????001?????1100011;
  parameter logic [31:0] C_ADD      = 32'b????????????????1001??????????10;
  parameter logic [31:0] C_ADDI     = 32'b????????????????000???????????01;
  parameter logic [31:0] C_ADDI16SP = 32'b????????????????011?00010?????01;
  parameter logic [31:0] C_ADDI4SPN = 32'b????????????????000???????????00;
  parameter logic [31:0] C_AND      = 32'b????????????????100011???11???01;
  parameter logic [31:0] C_ANDI     = 32'b????????????????100?10????????01;
  parameter logic [31:0] C_BEQZ     = 32'b????????????????110???????????01;
  parameter logic [31:0] C_BNEZ     = 32'b????????????????111???????????01;
  parameter logic [31:0] C_EBREAK   = 32'b????????????????1001000000000010;
  parameter logic [31:0] C_JALR     = 32'b????????????????1001?????0000010;
  parameter logic [31:0] C_JAL      = 32'b????????????????001???????????01;
  parameter logic [31:0] C_JR       = 32'b????????????????1000?????0000010;
  parameter logic [31:0] C_LI       = 32'b????????????????010???????????01;
  parameter logic [31:0] C_LUI      = 32'b????????????????011???????????01;
  parameter logic [31:0] C_LW       = 32'b????????????????010???????????00;
  parameter logic [31:0] C_LWSP     = 32'b????????????????010???????????10;
  parameter logic [31:0] C_MV       = 32'b????????????????1000??????????10;
  parameter logic [31:0] C_NOP      = 32'b????????????????000?00000?????01;
  parameter logic [31:0] C_OR       = 32'b????????????????100011???10???01;
  parameter logic [31:0] C_SUB      = 32'b????????????????100011???00???01;
  parameter logic [31:0] C_SW       = 32'b????????????????110???????????00;
  parameter logic [31:0] C_SWSP     = 32'b????????????????110???????????10;
  parameter logic [31:0] C_XOR      = 32'b????????????????100011???01???01;
  parameter logic [31:0] CSRRC      = 32'b?????????????????011?????1110011;
  parameter logic [31:0] CSRRCI     = 32'b?????????????????111?????1110011;
  parameter logic [31:0] CSRRS      = 32'b?????????????????010?????1110011;
  parameter logic [31:0] CSRRSI     = 32'b?????????????????110?????1110011;
  parameter logic [31:0] CSRRW      = 32'b?????????????????001?????1110011;
  parameter logic [31:0] CSRRWI     = 32'b?????????????????101?????1110011;
  parameter logic [31:0] DIV        = 32'b0000001??????????100?????0110011;
  parameter logic [31:0] DIVU       = 32'b0000001??????????101?????0110011;
  parameter logic [31:0] EBREAK     = 32'b00000000000100000000000001110011;
  parameter logic [31:0] ECALL      = 32'b00000000000000000000000001110011;
  parameter logic [31:0] FENCE      = 32'b?????????????????000?????0001111;
  parameter logic [31:0] JALR       = 32'b?????????????????000?????1100111;
  parameter logic [31:0] LB         = 32'b?????????????????000?????0000011;
  parameter logic [31:0] LBU        = 32'b?????????????????100?????0000011;
  parameter logic [31:0] LH         = 32'b?????????????????001?????0000011;
  parameter logic [31:0] LHU        = 32'b?????????????????101?????0000011;
  parameter logic [31:0] LUI        = 32'b?????????????????????????0110111;
  parameter logic [31:0] LW         = 32'b?????????????????010?????0000011;
  parameter logic [31:0] MRET       = 32'b00110000001000000000000001110011;
  parameter logic [31:0] MUL        = 32'b0000001??????????000?????0110011;
  parameter logic [31:0] MULH       = 32'b0000001??????????001?????0110011;
  parameter logic [31:0] MULHSU     = 32'b0000001??????????010?????0110011;
  parameter logic [31:0] MULHU      = 32'b0000001??????????011?????0110011;
  parameter logic [31:0] OR         = 32'b0000000??????????110?????0110011;
  parameter logic [31:0] ORI        = 32'b?????????????????110?????0010011;
  parameter logic [31:0] REM        = 32'b0000001??????????110?????0110011;
  parameter logic [31:0] REMU       = 32'b0000001??????????111?????0110011;
  parameter logic [31:0] SB         = 32'b?????????????????000?????0100011;
  parameter logic [31:0] SH         = 32'b?????????????????001?????0100011;
  parameter logic [31:0] SLL        = 32'b0000000??????????001?????0110011;
  parameter logic [31:0] SLLI       = 32'b0000000??????????001?????0010011;
  parameter logic [31:0] SLT        = 32'b0000000??????????010?????0110011;
  parameter logic [31:0] SLTI       = 32'b?????????????????010?????0010011;
  parameter logic [31:0] SLTIU      = 32'b?????????????????011?????0010011;
  parameter logic [31:0] SLTU       = 32'b0000000??????????011?????0110011;
  parameter logic [31:0] SRA        = 32'b0100000??????????101?????0110011;
  parameter logic [31:0] SRAI       = 32'b0100000??????????101?????0010011;
  parameter logic [31:0] SRL        = 32'b0000000??????????101?????0110011;
  parameter logic [31:0] SRLI       = 32'b0000000??????????101?????0010011;
  parameter logic [31:0] SUB        = 32'b0100000??????????000?????0110011;
  parameter logic [31:0] SW         = 32'b?????????????????010?????0100011;
  parameter logic [31:0] WFI        = 32'b00010000010100000000000001110011;
  parameter logic [31:0] XOR        = 32'b0000000??????????100?????0110011;
  parameter logic [31:0] XORI       = 32'b?????????????????100?????0010011;
  parameter logic [31:0] C_J        = 32'b????????????????101???????????01;
  parameter logic [31:0] JAL        = 32'b?????????????????????????1101111;
  parameter logic [31:0] C_ILLEGAL  = 32'b????????????????0000000000000000;
  parameter logic [31:0] C_SLLI     = 32'b????????????????000???????????10;
  parameter logic [31:0] C_SRAI     = 32'b????????????????100?01????????01;
  parameter logic [31:0] C_SRLI     = 32'b????????????????100?00????????01;
  parameter logic [31:0] FENCEI     = 32'b00000000000000000001000000001111;
  // verilog_format: on

  // verilog_format: off
  parameter logic [2:0] AluAddFunct3     = 3'b000;
  parameter logic [2:0] AluSubFunct3     = 3'b000;

  parameter logic [2:0] AluSllFunct3     = 3'b001;
  parameter logic [2:0] AluSltFunct3     = 3'b010;
  parameter logic [2:0] AluSltuFunct3    = 3'b011;
  parameter logic [2:0] AluXorFunct3     = 3'b100;

  parameter logic [2:0] AluSrlFunct3     = 3'b101;
  parameter logic [2:0] AluSraFunct3     = 3'b101;

  parameter logic [2:0] AluOrFunct3      = 3'b110;
  parameter logic [2:0] AluAndFunct3     = 3'b111;

  parameter logic [2:0] AluMulFunct3     = 3'b000;
  parameter logic [2:0] AluMulhFunct3    = 3'b001;
  parameter logic [2:0] AluMulhsuFunct3  = 3'b010;
  parameter logic [2:0] AluMulhuFunct3   = 3'b011;

  parameter logic [2:0] AluDivFunct3     = 3'b100;
  parameter logic [2:0] AluDivuFunct3    = 3'b101;
  parameter logic [2:0] AluRemFunct3     = 3'b110;
  parameter logic [2:0] AluRemuFunct3    = 3'b111;

  parameter logic [1:0] AluBasePrepend   = 2'b00;
  parameter logic [1:0] AluSubSraPrepend = 2'b01;
  parameter logic [1:0] AluMulPrepend    = 2'b11;
  // verilog_format: on

  // verilog_format: off
  parameter logic [4:0] ALU_ADD    = {{AluBasePrepend,   AluAddFunct3}};
  parameter logic [4:0] ALU_SUB    = {{AluSubSraPrepend, AluSubFunct3}};

  parameter logic [4:0] ALU_SLT    = {{AluBasePrepend,   AluSltFunct3}};
  parameter logic [4:0] ALU_SLTU   = {{AluBasePrepend,   AluSltuFunct3}};
  parameter logic [4:0] ALU_XOR    = {{AluBasePrepend,   AluXorFunct3}};
  parameter logic [4:0] ALU_OR     = {{AluBasePrepend,   AluOrFunct3}};
  parameter logic [4:0] ALU_AND    = {{AluBasePrepend,   AluAndFunct3}};
  parameter logic [4:0] ALU_SLL    = {{AluBasePrepend,   AluSllFunct3}};
  parameter logic [4:0] ALU_SRL    = {{AluBasePrepend,   AluSrlFunct3}};

  parameter logic [4:0] ALU_SRA    = {{AluSubSraPrepend, AluSraFunct3}};

  parameter logic [4:0] ALU_MUL    = {{AluMulPrepend,    AluMulFunct3}};
  parameter logic [4:0] ALU_MULH   = {{AluMulPrepend,    AluMulhFunct3}};
  parameter logic [4:0] ALU_MULHSU = {{AluMulPrepend,    AluMulhsuFunct3}};
  parameter logic [4:0] ALU_MULHU  = {{AluMulPrepend,    AluMulhuFunct3}};
  parameter logic [4:0] ALU_DIV    = {{AluMulPrepend,    AluDivFunct3}};
  parameter logic [4:0] ALU_DIVU   = {{AluMulPrepend,    AluDivuFunct3}};
  parameter logic [4:0] ALU_REM    = {{AluMulPrepend,    AluRemFunct3}};
  parameter logic [4:0] ALU_REMU   = {{AluMulPrepend,    AluRemuFunct3}};
  // verilog_format: on

  /*
   * Logic[3]: 0 -> Load, 1 -> Store
   * Logic[2]: 0 -> Signed, 1 -> Unsigned (LBU and LHU only)
   * Logic[1-0]: 00 -> Byte,  ?1 -> Half, 10 -> Word
   */

  // verilog_format: off
  parameter logic [3:0] LSU_LB  = 4'b0000;
  parameter logic [3:0] LSU_LH  = 4'b00?1;
  parameter logic [3:0] LSU_LW  = 4'b0010;
  parameter logic [3:0] LSU_LBU = 4'b0100;
  parameter logic [3:0] LSU_LHU = 4'b01?1;
  parameter logic [3:0] LSU_SB  = 4'b1000;
  parameter logic [3:0] LSU_SH  = 4'b10?1;
  parameter logic [3:0] LSU_SW  = 4'b1010;
  // verilog_format: on

  // verilog_format: off
  parameter logic [2:0] BR_BEQ  = 3'b000;
  parameter logic [2:0] BR_BGE  = 3'b101;
  parameter logic [2:0] BR_BGEU = 3'b111;
  parameter logic [2:0] BR_BNEZ = 3'b011;
  parameter logic [2:0] BR_BLT  = 3'b100;
  parameter logic [2:0] BR_BLTU = 3'b110;
  parameter logic [2:0] BR_BEQZ = 3'b010;
  parameter logic [2:0] BR_BNE  = 3'b001;
  // verilog_format: on

  // verilog_format: off
  parameter logic [1:0] FIXED  = 2'b00;
  parameter logic [1:0] INCR   = 2'b01;
  parameter logic [1:0] WRAP   = 2'b10;

  parameter logic [1:0] OKAY   = 2'b00;
  parameter logic [1:0] EXOKAY = 2'b01;
  parameter logic [1:0] SLVERR = 2'b10;
  parameter logic [1:0] DECERR = 2'b11;
  // verilog_format: on

  // Do not change these values.

  // verilog_format: off
  parameter int AddrW     = 32;
  parameter int DataW     = 32;
  parameter int RegCount  = 32;
  parameter int RegAddrW  = (RegCount > 1) ? $clog2(RegCount) : 0;
  parameter int AluOpW    = 5;
  parameter int LsuOpW    = 4;
  parameter int BranchOpW = 3;
  parameter int AxiIdW    = 2;
  // verilog_format: on

  // verilog_format: off
  parameter logic [31:0] Nop  = 32'h13;
  // verilog_format: on

endpackage
