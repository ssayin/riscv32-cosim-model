`ifndef DEC_DECODE_REF_MODEL_PKG
`define DEC_DECODE_REF_MODEL_PKG

package dec_decode_ref_model_pkg;

  import uvm_pkg::*;

  `include "uvm_macros.svh"

  import dec_decode_agent_pkg::*;

  `include "dec_decode_ref_model.sv"

endpackage : dec_decode_ref_model_pkg

`endif
