../../../../src/rtl/core/riscv_core.sv