// SPDX-FileCopyrightText: 2023 Serdar Sayın <https://serdarsayin.com>
//
// SPDX-License-Identifier: Apache-2.0

//=============================================================================
// Project  : src/tb/uvm_top
//
// File Name: top_tb.sv
//
// Author   : Name   : Serdar Sayın
//            Email  : serdarsayin@pm.me
//            Year   : 2023
//
// Version:   0.1
//
// Code created by Easier UVM Code Generator version 2017-01-19 on Thu Aug 10 23:43:50 2023
//=============================================================================
// Description: Testbench
//=============================================================================

module top_untimed_tb;

  timeunit      1ns;
  timeprecision 1ps;

  `include "uvm_macros.svh"

  import uvm_pkg::*;

  import top_test_pkg::*;
  import top_pkg::top_config;

  // Configuration object for top-level environment
  top_config top_env_config;

  // You can insert code here by setting tb_inc_inside_module in file tools/gen/common.tpl

  // You can remove the initial block below by setting tb_generate_run_test = no in file tools/gen/common.tpl

  initial
  begin
    // You can insert code here by setting tb_prepend_to_initial in file tools/gen/common.tpl

    // Create and populate top-level configuration object
    top_env_config = new("top_env_config");
    if ( !top_env_config.randomize() )
      `uvm_error("top_untimed_tb", "Failed to randomize top-level configuration object" )

    top_env_config.m_axi4master_config.vif = top_hdl_th.axi4master_bfm_0;

    uvm_config_db #(top_config)::set(null, "uvm_test_top", "config", top_env_config);
    uvm_config_db #(top_config)::set(null, "uvm_test_top.m_env", "config", top_env_config);

    // You can insert code here by setting tb_inc_before_run_test in file tools/gen/common.tpl

    run_test();
  end

endmodule

