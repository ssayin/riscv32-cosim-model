../../../../src/rtl/include/instr_defs.sv