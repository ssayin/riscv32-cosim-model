`ifndef DEC_DECODE_SEQ_LIST
`define DEC_DECODE_SEQ_LIST

package dec_decode_seq_list;

  import uvm_pkg::*;

  `include "uvm_macros.svh"

  import dec_decode_agent_pkg::*;
  import dec_decode_ref_model_pkg::*;
  import dec_decode_env_pkg::*;

  `include "dec_decode_basic_seq.sv"
  `include "dec_decode_instr_seq_from_file.sv"

endpackage : dec_decode_seq_list

`endif
