// SPDX-FileCopyrightText: 2023 Serdar Sayın <https://serdarsayin.com>
//
// SPDX-License-Identifier: Apache-2.0

package mem_stage_pkg;

  import uvm_pkg::*;

  `include "uvm_macros.svh"

  `include "mem_stage_agent.sv"
  `include "mem_stage_monitor.sv"
  `include "mem_stage_driver.sv"
  `include "mem_stage_sequencer.sv"
  `include "mem_stage_sequence.sv"

endpackage : mem_stage_pkg
