// SPDX-FileCopyrightText: 2023 Serdar Sayın <https://serdarsayin.com>
//
// SPDX-License-Identifier: Apache-2.0

//=============================================================================
// Project  : src/tb/uvm_top
//
// File Name: axi4master_sequencer.sv
//
// Author   : Name   : Serdar Sayın
//            Email  : serdarsayin@pm.me
//            Year   : 2023
//
// Version:   0.1
//
// Code created by Easier UVM Code Generator version 2017-01-19 on Thu Aug 10 23:12:34 2023
//=============================================================================
// Description: Sequencer for axi4master
//=============================================================================

`ifndef AXI4MASTER_SEQUENCER_SV
`define AXI4MASTER_SEQUENCER_SV

// Sequencer class is specialization of uvm_sequencer
typedef uvm_sequencer #(axi4_tx) axi4master_sequencer_t;


`endif // AXI4MASTER_SEQUENCER_SV

