// SPDX-FileCopyrightText: 2023 Serdar Sayın <https://serdarsayin.com>
//
// SPDX-License-Identifier: Apache-2.0

//=============================================================================
// Project  : src/tb/uvm_top
//
// File Name: axi4master_seq_lib.sv
//
// Author   : Name   : Serdar Sayın
//            Email  : serdarsayin@pm.me
//            Year   : 2023
//
// Version:   0.1
//
// Code created by Easier UVM Code Generator version 2017-01-19 on Thu Aug 10 23:12:34 2023
//=============================================================================
// Description: Sequence for agent axi4master
//=============================================================================

`ifndef AXI4MASTER_SEQ_LIB_SV
`define AXI4MASTER_SEQ_LIB_SV

class axi4master_default_seq extends uvm_sequence #(axi4_tx);

  `uvm_object_utils(axi4master_default_seq)

  axi4master_config  m_config;

  extern function new(string name = "");
  extern task body();

`ifndef UVM_POST_VERSION_1_1
  // Functions to support UVM 1.2 objection API in UVM 1.1
  extern function uvm_phase get_starting_phase();
  extern function void set_starting_phase(uvm_phase phase);
`endif

endclass : axi4master_default_seq


function axi4master_default_seq::new(string name = "");
  super.new(name);
endfunction : new


task axi4master_default_seq::body();
  `uvm_info(get_type_name(), "Default sequence starting", UVM_HIGH)

  req = axi4_tx::type_id::create("req");
  start_item(req); 
  if ( !req.randomize() )
    `uvm_error(get_type_name(), "Failed to randomize transaction")
  finish_item(req); 

  `uvm_info(get_type_name(), "Default sequence completed", UVM_HIGH)
endtask : body


`ifndef UVM_POST_VERSION_1_1
function uvm_phase axi4master_default_seq::get_starting_phase();
  return starting_phase;
endfunction: get_starting_phase


function void axi4master_default_seq::set_starting_phase(uvm_phase phase);
  starting_phase = phase;
endfunction: set_starting_phase
`endif


// Start of inlined include file src/tb/uvm_top/tb/include/my_axi4master_seq.sv
`ifndef MY_AXI4MASTER_SEQ_SV
`define MY_AXI4MASTER_SEQ_SV

class axi4master_hex_seq extends axi4master_default_seq;

  `uvm_object_utils(axi4master_hex_seq)

  function new(string name = "axi4master_hex_seq");
    super.new(name);
  endfunction : new

  task body();
    `uvm_info(get_type_name(), "axi4master_hex_seq sequence starting", UVM_HIGH)

    req = axi4_tx::type_id::create("req");

    start_item(req);

    assert (req.randomize() with {rid == 2'b00;});

    finish_item(req);

    `uvm_info(get_type_name(), "axi4master_hex_seq sequence completed", UVM_HIGH)
  endtask : body
endclass : axi4master_hex_seq

class axi4master_instr_feed_seq extends axi4master_default_seq;

  `uvm_object_utils(axi4master_instr_feed_seq)

  int          fd;
  logic [31:0] data[2];

  function new(string name = "axi4master_instr_feed_seq");
    super.new(name);
    fd = $fopen(`INSTR_SEQ_FILENAME, "r");
  endfunction : new

  task body();
    `uvm_info(get_type_name(), "axi4master_instr_feed_seq sequence starting", UVM_HIGH)


    for (int i = 0; i < `INSTR_SEQ_LINECOUNT / 2; ++i) begin
      req = axi4_tx::type_id::create("req");

      // TODO: fix endian
      for (int i = 0; i < 2; i++) begin
        $fscanf(fd, "%d", data[i]);
      end

      start_item(req);

      assert (req.randomize() with {rid == 2'b00;});
      for (int i = 0; i < 2; i++) begin
        // TODO: fix endian
        req.rdata[i] = data[i];
      end

      finish_item(req);
    end

    $fclose(fd);
    `uvm_info(get_type_name(), "axi4master_instr_feed_seq sequence completed", UVM_HIGH)
  endtask : body

endclass : axi4master_instr_feed_seq

`endif
// End of inlined include file

`endif // AXI4MASTER_SEQ_LIB_SV

