uvm_analysis_export #(riscv_core_tx) analysis_port = new("analysis_port", this);
axi4_logic m_axi4_logic = new();
