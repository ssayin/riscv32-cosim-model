
module platform (
	clk_clk,
	rst_n_reset_n);	

	input		clk_clk;
	input		rst_n_reset_n;
endmodule
