module riscv_decoder_j_no_rr (
  input  logic [15:0] instr,
  output logic        j
);
  always_comb begin
    casez (instr)
      16'b?????????1101111: j = 1;
      16'b?01???????????01: j = 1;
      default:              j = 0;
    endcase
  end

endmodule
