../../../../src/rtl/include/param_defs.sv