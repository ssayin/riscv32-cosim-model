import defs_pkg::*;
module ifu_br ();
endmodule
