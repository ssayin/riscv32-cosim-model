// platform.v

// Generated using ACDS version 22.1 917

`timescale 1 ps / 1 ps
module platform (
		input  wire  clk_clk,       //   clk.clk
		input  wire  rst_n_reset_n  // rst_n.reset_n
	);

	wire   [1:0] riscv_core_0_altera_axi4_master_1_awburst;                  // riscv_core_0:axi_awburst -> mm_interconnect_0:riscv_core_0_altera_axi4_master_1_awburst
	wire   [3:0] riscv_core_0_altera_axi4_master_1_arregion;                 // riscv_core_0:axi_arregion -> mm_interconnect_0:riscv_core_0_altera_axi4_master_1_arregion
	wire   [7:0] riscv_core_0_altera_axi4_master_1_arlen;                    // riscv_core_0:axi_arlen -> mm_interconnect_0:riscv_core_0_altera_axi4_master_1_arlen
	wire   [3:0] riscv_core_0_altera_axi4_master_1_arqos;                    // riscv_core_0:axi_arqos -> mm_interconnect_0:riscv_core_0_altera_axi4_master_1_arqos
	wire   [7:0] riscv_core_0_altera_axi4_master_1_wstrb;                    // riscv_core_0:axi_wstrb -> mm_interconnect_0:riscv_core_0_altera_axi4_master_1_wstrb
	wire         riscv_core_0_altera_axi4_master_1_wready;                   // mm_interconnect_0:riscv_core_0_altera_axi4_master_1_wready -> riscv_core_0:axi_wready
	wire         riscv_core_0_altera_axi4_master_1_rid;                      // mm_interconnect_0:riscv_core_0_altera_axi4_master_1_rid -> riscv_core_0:axi_rid
	wire         riscv_core_0_altera_axi4_master_1_rready;                   // riscv_core_0:axi_rready -> mm_interconnect_0:riscv_core_0_altera_axi4_master_1_rready
	wire   [7:0] riscv_core_0_altera_axi4_master_1_awlen;                    // riscv_core_0:axi_awlen -> mm_interconnect_0:riscv_core_0_altera_axi4_master_1_awlen
	wire   [3:0] riscv_core_0_altera_axi4_master_1_awqos;                    // riscv_core_0:axi_awqos -> mm_interconnect_0:riscv_core_0_altera_axi4_master_1_awqos
	wire   [3:0] riscv_core_0_altera_axi4_master_1_arcache;                  // riscv_core_0:axi_arcache -> mm_interconnect_0:riscv_core_0_altera_axi4_master_1_arcache
	wire         riscv_core_0_altera_axi4_master_1_wvalid;                   // riscv_core_0:axi_wvalid -> mm_interconnect_0:riscv_core_0_altera_axi4_master_1_wvalid
	wire  [31:0] riscv_core_0_altera_axi4_master_1_araddr;                   // riscv_core_0:axi_araddr -> mm_interconnect_0:riscv_core_0_altera_axi4_master_1_araddr
	wire   [2:0] riscv_core_0_altera_axi4_master_1_arprot;                   // riscv_core_0:axi_arprot -> mm_interconnect_0:riscv_core_0_altera_axi4_master_1_arprot
	wire   [2:0] riscv_core_0_altera_axi4_master_1_awprot;                   // riscv_core_0:axi_awprot -> mm_interconnect_0:riscv_core_0_altera_axi4_master_1_awprot
	wire  [63:0] riscv_core_0_altera_axi4_master_1_wdata;                    // riscv_core_0:axi_wdata -> mm_interconnect_0:riscv_core_0_altera_axi4_master_1_wdata
	wire         riscv_core_0_altera_axi4_master_1_arvalid;                  // riscv_core_0:axi_arvalid -> mm_interconnect_0:riscv_core_0_altera_axi4_master_1_arvalid
	wire   [3:0] riscv_core_0_altera_axi4_master_1_awcache;                  // riscv_core_0:axi_awcache -> mm_interconnect_0:riscv_core_0_altera_axi4_master_1_awcache
	wire         riscv_core_0_altera_axi4_master_1_arid;                     // riscv_core_0:axi_arid -> mm_interconnect_0:riscv_core_0_altera_axi4_master_1_arid
	wire         riscv_core_0_altera_axi4_master_1_arlock;                   // riscv_core_0:axi_arlock -> mm_interconnect_0:riscv_core_0_altera_axi4_master_1_arlock
	wire         riscv_core_0_altera_axi4_master_1_awlock;                   // riscv_core_0:axi_awlock -> mm_interconnect_0:riscv_core_0_altera_axi4_master_1_awlock
	wire  [31:0] riscv_core_0_altera_axi4_master_1_awaddr;                   // riscv_core_0:axi_awaddr -> mm_interconnect_0:riscv_core_0_altera_axi4_master_1_awaddr
	wire   [1:0] riscv_core_0_altera_axi4_master_1_bresp;                    // mm_interconnect_0:riscv_core_0_altera_axi4_master_1_bresp -> riscv_core_0:axi_bresp
	wire         riscv_core_0_altera_axi4_master_1_arready;                  // mm_interconnect_0:riscv_core_0_altera_axi4_master_1_arready -> riscv_core_0:axi_arready
	wire  [63:0] riscv_core_0_altera_axi4_master_1_rdata;                    // mm_interconnect_0:riscv_core_0_altera_axi4_master_1_rdata -> riscv_core_0:axi_rdata
	wire         riscv_core_0_altera_axi4_master_1_awready;                  // mm_interconnect_0:riscv_core_0_altera_axi4_master_1_awready -> riscv_core_0:axi_awready
	wire   [1:0] riscv_core_0_altera_axi4_master_1_arburst;                  // riscv_core_0:axi_arburst -> mm_interconnect_0:riscv_core_0_altera_axi4_master_1_arburst
	wire   [2:0] riscv_core_0_altera_axi4_master_1_arsize;                   // riscv_core_0:axi_arsize -> mm_interconnect_0:riscv_core_0_altera_axi4_master_1_arsize
	wire         riscv_core_0_altera_axi4_master_1_bready;                   // riscv_core_0:axi_bready -> mm_interconnect_0:riscv_core_0_altera_axi4_master_1_bready
	wire         riscv_core_0_altera_axi4_master_1_rlast;                    // mm_interconnect_0:riscv_core_0_altera_axi4_master_1_rlast -> riscv_core_0:axi_rlast
	wire         riscv_core_0_altera_axi4_master_1_wlast;                    // riscv_core_0:axi_wlast -> mm_interconnect_0:riscv_core_0_altera_axi4_master_1_wlast
	wire   [3:0] riscv_core_0_altera_axi4_master_1_awregion;                 // riscv_core_0:axi_awregion -> mm_interconnect_0:riscv_core_0_altera_axi4_master_1_awregion
	wire   [1:0] riscv_core_0_altera_axi4_master_1_rresp;                    // mm_interconnect_0:riscv_core_0_altera_axi4_master_1_rresp -> riscv_core_0:axi_rresp
	wire         riscv_core_0_altera_axi4_master_1_awid;                     // riscv_core_0:axi_awid -> mm_interconnect_0:riscv_core_0_altera_axi4_master_1_awid
	wire         riscv_core_0_altera_axi4_master_1_bid;                      // mm_interconnect_0:riscv_core_0_altera_axi4_master_1_bid -> riscv_core_0:axi_bid
	wire         riscv_core_0_altera_axi4_master_1_bvalid;                   // mm_interconnect_0:riscv_core_0_altera_axi4_master_1_bvalid -> riscv_core_0:axi_bvalid
	wire   [2:0] riscv_core_0_altera_axi4_master_1_awsize;                   // riscv_core_0:axi_awsize -> mm_interconnect_0:riscv_core_0_altera_axi4_master_1_awsize
	wire         riscv_core_0_altera_axi4_master_1_awvalid;                  // riscv_core_0:axi_awvalid -> mm_interconnect_0:riscv_core_0_altera_axi4_master_1_awvalid
	wire         riscv_core_0_altera_axi4_master_1_rvalid;                   // mm_interconnect_0:riscv_core_0_altera_axi4_master_1_rvalid -> riscv_core_0:axi_rvalid
	wire  [31:0] mm_interconnect_0_ssram_0_avalon_ssram_slave_readdata;      // ssram_0:avalon_ssram_slave_readdata -> mm_interconnect_0:ssram_0_avalon_ssram_slave_readdata
	wire         mm_interconnect_0_ssram_0_avalon_ssram_slave_waitrequest;   // ssram_0:avalon_ssram_slave_waitrequest -> mm_interconnect_0:ssram_0_avalon_ssram_slave_waitrequest
	wire         mm_interconnect_0_ssram_0_avalon_ssram_slave_debugaccess;   // mm_interconnect_0:ssram_0_avalon_ssram_slave_debugaccess -> ssram_0:avalon_ssram_slave_debugaccess
	wire  [19:0] mm_interconnect_0_ssram_0_avalon_ssram_slave_address;       // mm_interconnect_0:ssram_0_avalon_ssram_slave_address -> ssram_0:avalon_ssram_slave_address
	wire         mm_interconnect_0_ssram_0_avalon_ssram_slave_read;          // mm_interconnect_0:ssram_0_avalon_ssram_slave_read -> ssram_0:avalon_ssram_slave_read
	wire   [3:0] mm_interconnect_0_ssram_0_avalon_ssram_slave_byteenable;    // mm_interconnect_0:ssram_0_avalon_ssram_slave_byteenable -> ssram_0:avalon_ssram_slave_byteenable
	wire         mm_interconnect_0_ssram_0_avalon_ssram_slave_readdatavalid; // ssram_0:avalon_ssram_slave_readdatavalid -> mm_interconnect_0:ssram_0_avalon_ssram_slave_readdatavalid
	wire         mm_interconnect_0_ssram_0_avalon_ssram_slave_lock;          // mm_interconnect_0:ssram_0_avalon_ssram_slave_lock -> ssram_0:avalon_ssram_slave_lock
	wire         mm_interconnect_0_ssram_0_avalon_ssram_slave_write;         // mm_interconnect_0:ssram_0_avalon_ssram_slave_write -> ssram_0:avalon_ssram_slave_write
	wire  [31:0] mm_interconnect_0_ssram_0_avalon_ssram_slave_writedata;     // mm_interconnect_0:ssram_0_avalon_ssram_slave_writedata -> ssram_0:avalon_ssram_slave_writedata
	wire   [2:0] mm_interconnect_0_ssram_0_avalon_ssram_slave_burstcount;    // mm_interconnect_0:ssram_0_avalon_ssram_slave_burstcount -> ssram_0:avalon_ssram_slave_burstcount

	riscv_core riscv_core_0 (
		.axi_awid     (riscv_core_0_altera_axi4_master_1_awid),     // altera_axi4_master_1.awid
		.axi_awaddr   (riscv_core_0_altera_axi4_master_1_awaddr),   //                     .awaddr
		.axi_awlen    (riscv_core_0_altera_axi4_master_1_awlen),    //                     .awlen
		.axi_awsize   (riscv_core_0_altera_axi4_master_1_awsize),   //                     .awsize
		.axi_awburst  (riscv_core_0_altera_axi4_master_1_awburst),  //                     .awburst
		.axi_awlock   (riscv_core_0_altera_axi4_master_1_awlock),   //                     .awlock
		.axi_awcache  (riscv_core_0_altera_axi4_master_1_awcache),  //                     .awcache
		.axi_awprot   (riscv_core_0_altera_axi4_master_1_awprot),   //                     .awprot
		.axi_awvalid  (riscv_core_0_altera_axi4_master_1_awvalid),  //                     .awvalid
		.axi_awregion (riscv_core_0_altera_axi4_master_1_awregion), //                     .awregion
		.axi_awqos    (riscv_core_0_altera_axi4_master_1_awqos),    //                     .awqos
		.axi_awready  (riscv_core_0_altera_axi4_master_1_awready),  //                     .awready
		.axi_wdata    (riscv_core_0_altera_axi4_master_1_wdata),    //                     .wdata
		.axi_wstrb    (riscv_core_0_altera_axi4_master_1_wstrb),    //                     .wstrb
		.axi_wlast    (riscv_core_0_altera_axi4_master_1_wlast),    //                     .wlast
		.axi_wvalid   (riscv_core_0_altera_axi4_master_1_wvalid),   //                     .wvalid
		.axi_wready   (riscv_core_0_altera_axi4_master_1_wready),   //                     .wready
		.axi_bid      (riscv_core_0_altera_axi4_master_1_bid),      //                     .bid
		.axi_bresp    (riscv_core_0_altera_axi4_master_1_bresp),    //                     .bresp
		.axi_bvalid   (riscv_core_0_altera_axi4_master_1_bvalid),   //                     .bvalid
		.axi_bready   (riscv_core_0_altera_axi4_master_1_bready),   //                     .bready
		.axi_arid     (riscv_core_0_altera_axi4_master_1_arid),     //                     .arid
		.axi_araddr   (riscv_core_0_altera_axi4_master_1_araddr),   //                     .araddr
		.axi_arlen    (riscv_core_0_altera_axi4_master_1_arlen),    //                     .arlen
		.axi_arsize   (riscv_core_0_altera_axi4_master_1_arsize),   //                     .arsize
		.axi_arburst  (riscv_core_0_altera_axi4_master_1_arburst),  //                     .arburst
		.axi_arlock   (riscv_core_0_altera_axi4_master_1_arlock),   //                     .arlock
		.axi_arcache  (riscv_core_0_altera_axi4_master_1_arcache),  //                     .arcache
		.axi_arprot   (riscv_core_0_altera_axi4_master_1_arprot),   //                     .arprot
		.axi_arvalid  (riscv_core_0_altera_axi4_master_1_arvalid),  //                     .arvalid
		.axi_arqos    (riscv_core_0_altera_axi4_master_1_arqos),    //                     .arqos
		.axi_arregion (riscv_core_0_altera_axi4_master_1_arregion), //                     .arregion
		.axi_arready  (riscv_core_0_altera_axi4_master_1_arready),  //                     .arready
		.axi_rid      (riscv_core_0_altera_axi4_master_1_rid),      //                     .rid
		.axi_rdata    (riscv_core_0_altera_axi4_master_1_rdata),    //                     .rdata
		.axi_rresp    (riscv_core_0_altera_axi4_master_1_rresp),    //                     .rresp
		.axi_rlast    (riscv_core_0_altera_axi4_master_1_rlast),    //                     .rlast
		.axi_rvalid   (riscv_core_0_altera_axi4_master_1_rvalid),   //                     .rvalid
		.axi_rready   (riscv_core_0_altera_axi4_master_1_rready),   //                     .rready
		.clk          (clk_clk),                                    //                  clk.clk
		.rst_n        (rst_n_reset_n)                               //                  rst.reset_n
	);

	platform_ssram_0 ssram_0 (
		.clk_clk                          (clk_clk),                                                    //                clk.clk
		.reset_reset_n                    (rst_n_reset_n),                                              //              reset.reset_n
		.avalon_ssram_slave_address       (mm_interconnect_0_ssram_0_avalon_ssram_slave_address),       // avalon_ssram_slave.address
		.avalon_ssram_slave_burstcount    (mm_interconnect_0_ssram_0_avalon_ssram_slave_burstcount),    //                   .burstcount
		.avalon_ssram_slave_read          (mm_interconnect_0_ssram_0_avalon_ssram_slave_read),          //                   .read
		.avalon_ssram_slave_write         (mm_interconnect_0_ssram_0_avalon_ssram_slave_write),         //                   .write
		.avalon_ssram_slave_waitrequest   (mm_interconnect_0_ssram_0_avalon_ssram_slave_waitrequest),   //                   .waitrequest
		.avalon_ssram_slave_readdatavalid (mm_interconnect_0_ssram_0_avalon_ssram_slave_readdatavalid), //                   .readdatavalid
		.avalon_ssram_slave_byteenable    (mm_interconnect_0_ssram_0_avalon_ssram_slave_byteenable),    //                   .byteenable
		.avalon_ssram_slave_readdata      (mm_interconnect_0_ssram_0_avalon_ssram_slave_readdata),      //                   .readdata
		.avalon_ssram_slave_writedata     (mm_interconnect_0_ssram_0_avalon_ssram_slave_writedata),     //                   .writedata
		.avalon_ssram_slave_lock          (mm_interconnect_0_ssram_0_avalon_ssram_slave_lock),          //                   .lock
		.avalon_ssram_slave_debugaccess   (mm_interconnect_0_ssram_0_avalon_ssram_slave_debugaccess),   //                   .debugaccess
		.external_interface_ssram_be_n    (),                                                           // external_interface.ssram_be_n
		.external_interface_ssram_we_n    (),                                                           //                   .ssram_we_n
		.external_interface_fs_dq         (),                                                           //                   .fs_dq
		.external_interface_ssram_adsc_n  (),                                                           //                   .ssram_adsc_n
		.external_interface_ssram_oe_n    (),                                                           //                   .ssram_oe_n
		.external_interface_fs_addr       (),                                                           //                   .fs_addr
		.external_interface_ssram_cs_n    ()                                                            //                   .ssram_cs_n
	);

	platform_mm_interconnect_0 mm_interconnect_0 (
		.riscv_core_0_altera_axi4_master_1_awid       (riscv_core_0_altera_axi4_master_1_awid),                     //      riscv_core_0_altera_axi4_master_1.awid
		.riscv_core_0_altera_axi4_master_1_awaddr     (riscv_core_0_altera_axi4_master_1_awaddr),                   //                                       .awaddr
		.riscv_core_0_altera_axi4_master_1_awlen      (riscv_core_0_altera_axi4_master_1_awlen),                    //                                       .awlen
		.riscv_core_0_altera_axi4_master_1_awsize     (riscv_core_0_altera_axi4_master_1_awsize),                   //                                       .awsize
		.riscv_core_0_altera_axi4_master_1_awburst    (riscv_core_0_altera_axi4_master_1_awburst),                  //                                       .awburst
		.riscv_core_0_altera_axi4_master_1_awlock     (riscv_core_0_altera_axi4_master_1_awlock),                   //                                       .awlock
		.riscv_core_0_altera_axi4_master_1_awcache    (riscv_core_0_altera_axi4_master_1_awcache),                  //                                       .awcache
		.riscv_core_0_altera_axi4_master_1_awprot     (riscv_core_0_altera_axi4_master_1_awprot),                   //                                       .awprot
		.riscv_core_0_altera_axi4_master_1_awqos      (riscv_core_0_altera_axi4_master_1_awqos),                    //                                       .awqos
		.riscv_core_0_altera_axi4_master_1_awregion   (riscv_core_0_altera_axi4_master_1_awregion),                 //                                       .awregion
		.riscv_core_0_altera_axi4_master_1_awvalid    (riscv_core_0_altera_axi4_master_1_awvalid),                  //                                       .awvalid
		.riscv_core_0_altera_axi4_master_1_awready    (riscv_core_0_altera_axi4_master_1_awready),                  //                                       .awready
		.riscv_core_0_altera_axi4_master_1_wdata      (riscv_core_0_altera_axi4_master_1_wdata),                    //                                       .wdata
		.riscv_core_0_altera_axi4_master_1_wstrb      (riscv_core_0_altera_axi4_master_1_wstrb),                    //                                       .wstrb
		.riscv_core_0_altera_axi4_master_1_wlast      (riscv_core_0_altera_axi4_master_1_wlast),                    //                                       .wlast
		.riscv_core_0_altera_axi4_master_1_wvalid     (riscv_core_0_altera_axi4_master_1_wvalid),                   //                                       .wvalid
		.riscv_core_0_altera_axi4_master_1_wready     (riscv_core_0_altera_axi4_master_1_wready),                   //                                       .wready
		.riscv_core_0_altera_axi4_master_1_bid        (riscv_core_0_altera_axi4_master_1_bid),                      //                                       .bid
		.riscv_core_0_altera_axi4_master_1_bresp      (riscv_core_0_altera_axi4_master_1_bresp),                    //                                       .bresp
		.riscv_core_0_altera_axi4_master_1_bvalid     (riscv_core_0_altera_axi4_master_1_bvalid),                   //                                       .bvalid
		.riscv_core_0_altera_axi4_master_1_bready     (riscv_core_0_altera_axi4_master_1_bready),                   //                                       .bready
		.riscv_core_0_altera_axi4_master_1_arid       (riscv_core_0_altera_axi4_master_1_arid),                     //                                       .arid
		.riscv_core_0_altera_axi4_master_1_araddr     (riscv_core_0_altera_axi4_master_1_araddr),                   //                                       .araddr
		.riscv_core_0_altera_axi4_master_1_arlen      (riscv_core_0_altera_axi4_master_1_arlen),                    //                                       .arlen
		.riscv_core_0_altera_axi4_master_1_arsize     (riscv_core_0_altera_axi4_master_1_arsize),                   //                                       .arsize
		.riscv_core_0_altera_axi4_master_1_arburst    (riscv_core_0_altera_axi4_master_1_arburst),                  //                                       .arburst
		.riscv_core_0_altera_axi4_master_1_arlock     (riscv_core_0_altera_axi4_master_1_arlock),                   //                                       .arlock
		.riscv_core_0_altera_axi4_master_1_arcache    (riscv_core_0_altera_axi4_master_1_arcache),                  //                                       .arcache
		.riscv_core_0_altera_axi4_master_1_arprot     (riscv_core_0_altera_axi4_master_1_arprot),                   //                                       .arprot
		.riscv_core_0_altera_axi4_master_1_arqos      (riscv_core_0_altera_axi4_master_1_arqos),                    //                                       .arqos
		.riscv_core_0_altera_axi4_master_1_arregion   (riscv_core_0_altera_axi4_master_1_arregion),                 //                                       .arregion
		.riscv_core_0_altera_axi4_master_1_arvalid    (riscv_core_0_altera_axi4_master_1_arvalid),                  //                                       .arvalid
		.riscv_core_0_altera_axi4_master_1_arready    (riscv_core_0_altera_axi4_master_1_arready),                  //                                       .arready
		.riscv_core_0_altera_axi4_master_1_rid        (riscv_core_0_altera_axi4_master_1_rid),                      //                                       .rid
		.riscv_core_0_altera_axi4_master_1_rdata      (riscv_core_0_altera_axi4_master_1_rdata),                    //                                       .rdata
		.riscv_core_0_altera_axi4_master_1_rresp      (riscv_core_0_altera_axi4_master_1_rresp),                    //                                       .rresp
		.riscv_core_0_altera_axi4_master_1_rlast      (riscv_core_0_altera_axi4_master_1_rlast),                    //                                       .rlast
		.riscv_core_0_altera_axi4_master_1_rvalid     (riscv_core_0_altera_axi4_master_1_rvalid),                   //                                       .rvalid
		.riscv_core_0_altera_axi4_master_1_rready     (riscv_core_0_altera_axi4_master_1_rready),                   //                                       .rready
		.clk_0_clk_clk                                (clk_clk),                                                    //                              clk_0_clk.clk
		.riscv_core_0_rst_reset_bridge_in_reset_reset (~rst_n_reset_n),                                             // riscv_core_0_rst_reset_bridge_in_reset.reset
		.ssram_0_reset_reset_bridge_in_reset_reset    (~rst_n_reset_n),                                             //    ssram_0_reset_reset_bridge_in_reset.reset
		.ssram_0_avalon_ssram_slave_address           (mm_interconnect_0_ssram_0_avalon_ssram_slave_address),       //             ssram_0_avalon_ssram_slave.address
		.ssram_0_avalon_ssram_slave_write             (mm_interconnect_0_ssram_0_avalon_ssram_slave_write),         //                                       .write
		.ssram_0_avalon_ssram_slave_read              (mm_interconnect_0_ssram_0_avalon_ssram_slave_read),          //                                       .read
		.ssram_0_avalon_ssram_slave_readdata          (mm_interconnect_0_ssram_0_avalon_ssram_slave_readdata),      //                                       .readdata
		.ssram_0_avalon_ssram_slave_writedata         (mm_interconnect_0_ssram_0_avalon_ssram_slave_writedata),     //                                       .writedata
		.ssram_0_avalon_ssram_slave_burstcount        (mm_interconnect_0_ssram_0_avalon_ssram_slave_burstcount),    //                                       .burstcount
		.ssram_0_avalon_ssram_slave_byteenable        (mm_interconnect_0_ssram_0_avalon_ssram_slave_byteenable),    //                                       .byteenable
		.ssram_0_avalon_ssram_slave_readdatavalid     (mm_interconnect_0_ssram_0_avalon_ssram_slave_readdatavalid), //                                       .readdatavalid
		.ssram_0_avalon_ssram_slave_waitrequest       (mm_interconnect_0_ssram_0_avalon_ssram_slave_waitrequest),   //                                       .waitrequest
		.ssram_0_avalon_ssram_slave_lock              (mm_interconnect_0_ssram_0_avalon_ssram_slave_lock),          //                                       .lock
		.ssram_0_avalon_ssram_slave_debugaccess       (mm_interconnect_0_ssram_0_avalon_ssram_slave_debugaccess)    //                                       .debugaccess
	);

endmodule
