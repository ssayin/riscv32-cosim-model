// TODO: what are trade-off btw. decompress expansion
// VS decode right justified w/ comp switch?

module ifu_aln ();

endmodule
