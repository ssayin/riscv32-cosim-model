// SPDX-FileCopyrightText: 2023 Serdar Sayın <https://serdarsayin.com>
//
// SPDX-License-Identifier: Apache-2.0

package ex_stage_pkg;

  import uvm_pkg::*;

  `include "uvm_macros.svh"

  `include "ex_stage_agent.sv"
  `include "ex_stage_monitor.sv"
  `include "ex_stage_driver.sv"
  `include "ex_stage_sequencer.sv"
  `include "ex_stage_sequence.sv"

endpackage : ex_stage_pkg
