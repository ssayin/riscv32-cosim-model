// SPDX-FileCopyrightText: 2023 Serdar Sayın <https://serdarsayin.com>
//
// SPDX-License-Identifier: Apache-2.0

//=============================================================================
// Project  : ../tb/uvm_top
//
// File Name: riscv_core_driver.sv
//
// Author   : Name   : Serdar Sayın
//            Email  : serdarsayin@pm.me
//            Year   : 2023
//
// Version:   0.1
//
// Code created by Easier UVM Code Generator version 2017-01-19 on Sat Jul 15 22:09:49 2023
//=============================================================================
// Description: Driver for riscv_core
//=============================================================================

`ifndef RISCV_CORE_DRIVER_SV
`define RISCV_CORE_DRIVER_SV

// You can insert code here by setting driver_inc_before_class in file riscv_core.tpl

class riscv_core_driver extends uvm_driver #(riscv_core_tx);

  `uvm_component_utils(riscv_core_driver)

  virtual riscv_core_if vif;

  riscv_core_config     m_config;

  extern function new(string name, uvm_component parent);

  // Methods run_phase and do_drive generated by setting driver_inc in file riscv_core.tpl
  extern task run_phase(uvm_phase phase);
  extern task do_drive();

  // You can insert code here by setting driver_inc_inside_class in file riscv_core.tpl

endclass : riscv_core_driver 


function riscv_core_driver::new(string name, uvm_component parent);
  super.new(name, parent);
endfunction : new


task riscv_core_driver::run_phase(uvm_phase phase);
  `uvm_info(get_type_name(), "run_phase", UVM_HIGH)

  forever
  begin
    seq_item_port.get_next_item(req);
      `uvm_info(get_type_name(), {"req item\n",req.sprint}, UVM_HIGH)
    do_drive();
    seq_item_port.item_done();
  end
endtask : run_phase


// Start of inlined include file ../tb/uvm_top/tb/include/riscv_core_do_drive.sv
task riscv_core_driver::do_drive();
  vif.mem_data_in[0] = req.mem_data_in[0];
  vif.mem_data_in[1] = req.mem_data_in[1];
  vif.mem_ready      = req.mem_ready;
  vif.irq_external   = req.irq_external;
  vif.irq_timer      = req.irq_timer;
  vif.irq_software   = req.irq_software;
  @(posedge vif.clk);
endtask
// End of inlined include file

// You can insert code here by setting driver_inc_after_class in file riscv_core.tpl

`endif // RISCV_CORE_DRIVER_SV

